TOOL:	xrun	23.09-s001: Started on Jan 16, 2026 at 08:57:11 EST
xrun: 23.09-s001: (c) Copyright 1995-2023 Cadence Design Systems, Inc.
	Top level design units:
		$unit_0x24a58354
		testbench
Loading snapshot worklib.testbench:sv .................... Done
SVSEED default: 1
xcelium> source /xcelium23.09/tools/xcelium/files/xmsimrc
xcelium> run
 GENERATOR CLASS DATA 
time =0,clk=0,rst=1,d=1,q=0
 DRIVER CLASS DATA 
time =5,clk=1,rst=1,d=1,q=0
 MONITOR CLASS DATA 
time =6,clk=1,rst=1,d=0,q=0
 SCOREBOARD CLASS DATA 
time =6,clk=1,rst=1,d=0,q=0
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =6,clk=1,rst=1,d=1,q=0
 DRIVER CLASS DATA 
time =15,clk=1,rst=0,d=1,q=0
 MONITOR CLASS DATA 
time =16,clk=1,rst=0,d=1,q=1
 SCOREBOARD CLASS DATA 
time =16,clk=1,rst=0,d=1,q=1
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =16,clk=1,rst=0,d=1,q=0
 DRIVER CLASS DATA 
time =25,clk=1,rst=0,d=1,q=0
 MONITOR CLASS DATA 
time =26,clk=1,rst=0,d=1,q=1
 SCOREBOARD CLASS DATA 
time =26,clk=1,rst=0,d=1,q=1
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =26,clk=1,rst=0,d=1,q=0
 DRIVER CLASS DATA 
time =35,clk=1,rst=0,d=1,q=0
 MONITOR CLASS DATA 
time =36,clk=1,rst=0,d=1,q=1
 SCOREBOARD CLASS DATA 
time =36,clk=1,rst=0,d=1,q=1
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =36,clk=1,rst=0,d=0,q=0
 DRIVER CLASS DATA 
time =45,clk=1,rst=0,d=0,q=0
 MONITOR CLASS DATA 
time =46,clk=1,rst=0,d=1,q=1
 SCOREBOARD CLASS DATA 
time =46,clk=1,rst=0,d=1,q=1
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =46,clk=1,rst=0,d=1,q=0
 DRIVER CLASS DATA 
time =55,clk=1,rst=0,d=1,q=0
 MONITOR CLASS DATA 
time =56,clk=1,rst=0,d=0,q=0
 SCOREBOARD CLASS DATA 
time =56,clk=1,rst=0,d=0,q=0
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =56,clk=1,rst=0,d=0,q=0
 DRIVER CLASS DATA 
time =65,clk=1,rst=0,d=0,q=0
 MONITOR CLASS DATA 
time =66,clk=1,rst=0,d=1,q=1
 SCOREBOARD CLASS DATA 
time =66,clk=1,rst=0,d=1,q=1
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =66,clk=1,rst=0,d=1,q=0
 DRIVER CLASS DATA 
time =75,clk=1,rst=0,d=1,q=0
 MONITOR CLASS DATA 
time =76,clk=1,rst=0,d=0,q=0
 SCOREBOARD CLASS DATA 
time =76,clk=1,rst=0,d=0,q=0
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =76,clk=1,rst=0,d=0,q=0
 DRIVER CLASS DATA 
time =85,clk=1,rst=0,d=0,q=0
 MONITOR CLASS DATA 
time =86,clk=1,rst=0,d=1,q=1
 SCOREBOARD CLASS DATA 
time =86,clk=1,rst=0,d=1,q=1
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =86,clk=1,rst=0,d=1,q=0
 DRIVER CLASS DATA 
time =95,clk=1,rst=0,d=1,q=0
 MONITOR CLASS DATA 
time =96,clk=1,rst=0,d=0,q=0
 SCOREBOARD CLASS DATA 
time =96,clk=1,rst=0,d=0,q=0
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =96,clk=1,rst=0,d=0,q=0
 DRIVER CLASS DATA 
time =105,clk=1,rst=0,d=0,q=0
 MONITOR CLASS DATA 
time =106,clk=1,rst=0,d=1,q=1
 SCOREBOARD CLASS DATA 
time =106,clk=1,rst=0,d=1,q=1
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =106,clk=1,rst=0,d=0,q=0
 DRIVER CLASS DATA 
time =115,clk=1,rst=0,d=0,q=0
 MONITOR CLASS DATA 
time =116,clk=1,rst=0,d=0,q=0
 SCOREBOARD CLASS DATA 
time =116,clk=1,rst=0,d=0,q=0
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =116,clk=1,rst=0,d=1,q=0
 DRIVER CLASS DATA 
time =125,clk=1,rst=0,d=1,q=0
 MONITOR CLASS DATA 
time =126,clk=1,rst=0,d=0,q=0
 SCOREBOARD CLASS DATA 
time =126,clk=1,rst=0,d=0,q=0
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =126,clk=1,rst=0,d=0,q=0
 DRIVER CLASS DATA 
time =135,clk=1,rst=0,d=0,q=0
 MONITOR CLASS DATA 
time =136,clk=1,rst=0,d=1,q=1
 SCOREBOARD CLASS DATA 
time =136,clk=1,rst=0,d=1,q=1
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =136,clk=1,rst=0,d=0,q=0
 DRIVER CLASS DATA 
time =145,clk=1,rst=0,d=0,q=0
 MONITOR CLASS DATA 
time =146,clk=1,rst=0,d=0,q=0
 SCOREBOARD CLASS DATA 
time =146,clk=1,rst=0,d=0,q=0
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =146,clk=1,rst=0,d=1,q=0
 DRIVER CLASS DATA 
time =155,clk=1,rst=0,d=1,q=0
 MONITOR CLASS DATA 
time =156,clk=1,rst=0,d=0,q=0
 SCOREBOARD CLASS DATA 
time =156,clk=1,rst=0,d=0,q=0
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =156,clk=1,rst=0,d=1,q=0
 DRIVER CLASS DATA 
time =165,clk=1,rst=0,d=1,q=0
 MONITOR CLASS DATA 
time =166,clk=1,rst=0,d=1,q=1
 SCOREBOARD CLASS DATA 
time =166,clk=1,rst=0,d=1,q=1
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =166,clk=1,rst=0,d=0,q=0
 DRIVER CLASS DATA 
time =175,clk=1,rst=0,d=0,q=0
 MONITOR CLASS DATA 
time =176,clk=1,rst=0,d=1,q=1
 SCOREBOARD CLASS DATA 
time =176,clk=1,rst=0,d=1,q=1
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =176,clk=1,rst=0,d=1,q=0
 DRIVER CLASS DATA 
time =185,clk=1,rst=0,d=1,q=0
 MONITOR CLASS DATA 
time =186,clk=1,rst=0,d=0,q=0
 SCOREBOARD CLASS DATA 
time =186,clk=1,rst=0,d=0,q=0
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =186,clk=1,rst=0,d=1,q=0
 DRIVER CLASS DATA 
time =195,clk=1,rst=0,d=1,q=0
 MONITOR CLASS DATA 
time =196,clk=1,rst=0,d=1,q=1
 SCOREBOARD CLASS DATA 
time =196,clk=1,rst=0,d=1,q=1
		PASS		
-----------------------------------------------		
Simulation complete via implicit call to $finish(1) at time 196 NS + 1
./test.sv:3 program test(intf vintf);
xcelium> exit
TOOL:	xrun	23.09-s001: Exiting on Jan 16, 2026 at 08:57:12 EST  (total: 00:00:01)
Done
